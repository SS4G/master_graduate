module PoolAddrGen(

);

endmodule