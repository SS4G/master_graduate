module Dense1_layer(
    
);

endmodule