module CNN_TopDesign(

);

Conv2D_1 conv2d_1_inst(
    clk,
    rst_n,
    enable,
    
    img_data_wr,
    img_data_in,
    
    pool_1_out_00,
    pool_1_out_01,
    pool_1_out_02,
    pool_1_out_03,
    pool_1_out_04,
    pool_1_out_05,
     
    pool_1_out_en
);


endmodule